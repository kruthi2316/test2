module sum(a,b,s);

input a, b;
output s;

assign s=a+b;
kruthi is a  cute piggy 

endmodule