module sum(a,b,s);

input a, b;
output s;

assign s=a+b;
kruthi is a  cute_test_1 piggy 

endmodule